module trig_chain (
    input           CLK1,
    input           CLK2,
    input           CLK3,
    input [3:0]     IDATA,
    output [3:0]    ODATA
);


    
endmodule